library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity CharRam is

    port (
        clka  : in  std_logic;
        wea   : in  std_logic;
        addra : in  std_logic_vector(10 downto 0);
        dina  : in  std_logic_vector(7 downto 0);
        douta : out std_logic_vector(7 downto 0);
        clkb  : in  std_logic;
        web   : in  std_logic;
        addrb : in  std_logic_vector(10 downto 0);
        dinb  : in  std_logic_vector(7 downto 0);
        doutb : out std_logic_vector(7 downto 0)
        );
end CharRam;

architecture BEHAVIORAL of CharRam is

-- Shared memory
    type ram_type is array (0 to 2047) of std_logic_vector (7 downto 0);
    shared variable RAM : ram_type := (
        x"00", x"00", x"38", x"44", x"04", x"34", x"4c", x"4c", x"38", x"00", x"00", x"00", x"00", x"1C", x"22", x"02",
        x"00", x"00", x"10", x"28", x"44", x"44", x"7c", x"44", x"44", x"00", x"00", x"00", x"1A", x"2A", x"2A", x"1C",
        x"00", x"00", x"78", x"24", x"24", x"38", x"24", x"24", x"78", x"00", x"00", x"00", x"00", x"08", x"14", x"22",
        x"00", x"00", x"38", x"44", x"40", x"40", x"40", x"44", x"38", x"00", x"00", x"00", x"22", x"3E", x"22", x"22",
        x"00", x"00", x"78", x"24", x"24", x"24", x"24", x"24", x"78", x"00", x"00", x"00", x"00", x"3C", x"12", x"12",
        x"00", x"00", x"7c", x"40", x"40", x"70", x"40", x"40", x"7c", x"00", x"00", x"00", x"1C", x"12", x"12", x"3C",
        x"00", x"00", x"7c", x"40", x"40", x"70", x"40", x"40", x"40", x"00", x"00", x"00", x"00", x"1C", x"22", x"20",
        x"00", x"00", x"38", x"44", x"40", x"40", x"4c", x"44", x"38", x"00", x"00", x"00", x"20", x"20", x"22", x"1C",
        x"00", x"00", x"44", x"44", x"44", x"7c", x"44", x"44", x"44", x"00", x"00", x"00", x"00", x"3C", x"12", x"12",
        x"00", x"00", x"38", x"10", x"10", x"10", x"10", x"10", x"38", x"00", x"00", x"00", x"12", x"12", x"12", x"3C",
        x"00", x"00", x"04", x"04", x"04", x"04", x"04", x"44", x"38", x"00", x"00", x"00", x"00", x"3E", x"20", x"20",
        x"00", x"00", x"44", x"48", x"50", x"60", x"50", x"48", x"44", x"00", x"00", x"00", x"38", x"20", x"20", x"3E",
        x"00", x"00", x"40", x"40", x"40", x"40", x"40", x"40", x"7c", x"00", x"00", x"00", x"00", x"3E", x"20", x"20",
        x"00", x"00", x"44", x"6c", x"54", x"54", x"44", x"44", x"44", x"00", x"00", x"00", x"38", x"20", x"20", x"20",
        x"00", x"00", x"44", x"44", x"64", x"54", x"4c", x"44", x"44", x"00", x"00", x"00", x"00", x"1E", x"20", x"20",
        x"00", x"00", x"38", x"44", x"44", x"44", x"44", x"44", x"38", x"00", x"00", x"00", x"26", x"22", x"22", x"1E",
        x"00", x"00", x"78", x"44", x"44", x"78", x"40", x"40", x"40", x"00", x"00", x"00", x"00", x"22", x"22", x"22",
        x"00", x"00", x"38", x"44", x"44", x"44", x"54", x"48", x"34", x"00", x"00", x"00", x"3E", x"22", x"22", x"22",
        x"00", x"00", x"78", x"44", x"44", x"78", x"50", x"48", x"44", x"00", x"00", x"00", x"00", x"1C", x"08", x"08",
        x"00", x"00", x"38", x"44", x"40", x"38", x"04", x"44", x"38", x"00", x"00", x"00", x"08", x"08", x"08", x"1C",
        x"00", x"00", x"7c", x"10", x"10", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", x"02", x"02", x"02",
        x"00", x"00", x"44", x"44", x"44", x"44", x"44", x"44", x"38", x"00", x"00", x"00", x"02", x"22", x"22", x"1C",
        x"00", x"00", x"44", x"44", x"44", x"28", x"28", x"10", x"10", x"00", x"00", x"00", x"00", x"22", x"24", x"28",
        x"00", x"00", x"44", x"44", x"44", x"44", x"54", x"6c", x"44", x"00", x"00", x"00", x"30", x"28", x"24", x"22",
        x"00", x"00", x"44", x"44", x"28", x"10", x"28", x"44", x"44", x"00", x"00", x"00", x"00", x"20", x"20", x"20",
        x"00", x"00", x"44", x"44", x"28", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"20", x"20", x"20", x"3E",
        x"00", x"00", x"7c", x"04", x"08", x"10", x"20", x"40", x"7c", x"00", x"00", x"00", x"00", x"22", x"36", x"2A",
        x"00", x"00", x"38", x"20", x"20", x"20", x"20", x"20", x"38", x"00", x"00", x"00", x"2A", x"22", x"22", x"22",
        x"00", x"00", x"00", x"40", x"20", x"10", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"22", x"32", x"2A",
        x"00", x"00", x"38", x"08", x"08", x"08", x"08", x"08", x"38", x"00", x"00", x"00", x"26", x"22", x"22", x"22",
        x"00", x"00", x"10", x"38", x"54", x"10", x"10", x"10", x"10", x"00", x"00", x"00", x"00", x"3E", x"22", x"22",
        x"00", x"00", x"00", x"10", x"20", x"7c", x"20", x"10", x"00", x"00", x"00", x"00", x"22", x"22", x"22", x"3E",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3C", x"22", x"22",
        x"00", x"00", x"10", x"10", x"10", x"10", x"10", x"00", x"10", x"00", x"00", x"00", x"3C", x"20", x"20", x"20",
        x"00", x"00", x"28", x"28", x"28", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"22", x"22",
        x"00", x"00", x"28", x"28", x"7c", x"28", x"7c", x"28", x"28", x"00", x"00", x"00", x"22", x"2A", x"24", x"1A",
        x"00", x"00", x"10", x"3c", x"50", x"38", x"14", x"78", x"10", x"00", x"00", x"00", x"00", x"3C", x"22", x"22",
        x"00", x"00", x"60", x"64", x"08", x"10", x"20", x"4c", x"0c", x"00", x"00", x"00", x"3C", x"28", x"24", x"22",
        x"00", x"00", x"20", x"50", x"50", x"20", x"54", x"48", x"34", x"00", x"00", x"00", x"00", x"1C", x"22", x"10",
        x"00", x"00", x"10", x"10", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"04", x"22", x"1C",
        x"00", x"00", x"08", x"10", x"20", x"20", x"20", x"10", x"08", x"00", x"00", x"00", x"00", x"3E", x"08", x"08",
        x"00", x"00", x"20", x"10", x"08", x"08", x"08", x"10", x"20", x"00", x"00", x"00", x"08", x"08", x"08", x"08",
        x"00", x"00", x"00", x"10", x"54", x"38", x"38", x"54", x"10", x"00", x"00", x"00", x"00", x"22", x"22", x"22",
        x"00", x"00", x"00", x"10", x"10", x"7c", x"10", x"10", x"00", x"00", x"00", x"00", x"22", x"22", x"22", x"1C",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"20", x"40", x"00", x"00", x"00", x"22", x"22", x"22",
        x"00", x"00", x"00", x"00", x"00", x"7c", x"00", x"00", x"00", x"00", x"00", x"00", x"14", x"14", x"08", x"08",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"10", x"00", x"00", x"00", x"00", x"22", x"22", x"22",
        x"00", x"00", x"00", x"04", x"08", x"10", x"20", x"40", x"00", x"00", x"00", x"00", x"2A", x"2A", x"36", x"22",
        x"00", x"00", x"38", x"44", x"4c", x"54", x"64", x"44", x"38", x"00", x"00", x"00", x"00", x"22", x"22", x"14",
        x"00", x"00", x"10", x"30", x"10", x"10", x"10", x"10", x"38", x"00", x"00", x"00", x"08", x"14", x"22", x"22",
        x"00", x"00", x"38", x"44", x"04", x"38", x"40", x"40", x"7c", x"00", x"00", x"00", x"00", x"22", x"22", x"14",
        x"00", x"00", x"38", x"44", x"04", x"08", x"04", x"44", x"38", x"00", x"00", x"00", x"08", x"08", x"08", x"08",
        x"00", x"00", x"08", x"18", x"28", x"48", x"7c", x"08", x"08", x"00", x"00", x"00", x"00", x"3E", x"02", x"04",
        x"00", x"00", x"7c", x"40", x"78", x"04", x"04", x"44", x"38", x"00", x"00", x"00", x"08", x"10", x"20", x"3E",
        x"00", x"00", x"38", x"40", x"40", x"78", x"44", x"44", x"38", x"00", x"00", x"00", x"00", x"38", x"20", x"20",
        x"00", x"00", x"7c", x"04", x"08", x"10", x"20", x"40", x"40", x"00", x"00", x"00", x"20", x"20", x"20", x"38",
        x"00", x"00", x"38", x"44", x"44", x"38", x"44", x"44", x"38", x"00", x"00", x"00", x"00", x"20", x"20", x"10",
        x"00", x"00", x"38", x"44", x"44", x"3c", x"04", x"04", x"38", x"00", x"00", x"00", x"08", x"04", x"02", x"02",
        x"00", x"00", x"00", x"00", x"10", x"00", x"00", x"10", x"00", x"00", x"00", x"00", x"00", x"0E", x"02", x"02",
        x"00", x"00", x"00", x"00", x"10", x"00", x"00", x"10", x"10", x"20", x"00", x"00", x"02", x"02", x"02", x"0E",
        x"00", x"00", x"08", x"10", x"20", x"40", x"20", x"10", x"08", x"00", x"00", x"00", x"00", x"08", x"1C", x"2A",
        x"00", x"00", x"00", x"00", x"7c", x"00", x"7c", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"08", x"08",
        x"00", x"00", x"20", x"10", x"08", x"04", x"08", x"10", x"20", x"00", x"00", x"00", x"00", x"00", x"08", x"10",
        x"00", x"00", x"38", x"44", x"04", x"08", x"10", x"00", x"10", x"00", x"00", x"00", x"3E", x"10", x"08", x"00",
        x"00", x"00", x"10", x"28", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"38", x"04", x"3c", x"44", x"3c", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"40", x"40", x"58", x"64", x"44", x"64", x"58", x"00", x"00", x"00", x"00", x"08", x"08", x"08",
        x"00", x"00", x"00", x"00", x"38", x"44", x"40", x"44", x"38", x"00", x"00", x"00", x"08", x"08", x"00", x"08",
        x"00", x"00", x"04", x"04", x"34", x"4c", x"44", x"4c", x"34", x"00", x"00", x"00", x"00", x"14", x"14", x"14",
        x"00", x"00", x"00", x"00", x"38", x"44", x"7c", x"40", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"08", x"14", x"10", x"38", x"10", x"10", x"10", x"00", x"00", x"00", x"00", x"14", x"14", x"36",
        x"00", x"00", x"00", x"00", x"34", x"4c", x"44", x"4c", x"34", x"04", x"38", x"00", x"00", x"36", x"14", x"14",
        x"00", x"00", x"40", x"40", x"58", x"64", x"44", x"44", x"44", x"00", x"00", x"00", x"00", x"08", x"1E", x"20",
        x"00", x"00", x"10", x"00", x"30", x"10", x"10", x"10", x"38", x"00", x"00", x"00", x"1C", x"02", x"3C", x"08",
        x"00", x"00", x"04", x"00", x"04", x"04", x"04", x"04", x"44", x"38", x"00", x"00", x"00", x"32", x"32", x"04",
        x"00", x"00", x"40", x"40", x"48", x"50", x"60", x"50", x"48", x"00", x"00", x"00", x"08", x"10", x"26", x"26",
        x"00", x"00", x"30", x"10", x"10", x"10", x"10", x"10", x"38", x"00", x"00", x"00", x"00", x"10", x"28", x"28",
        x"00", x"00", x"00", x"00", x"78", x"54", x"54", x"54", x"54", x"00", x"00", x"00", x"10", x"2A", x"24", x"1A",
        x"00", x"00", x"00", x"00", x"58", x"64", x"44", x"44", x"44", x"00", x"00", x"00", x"00", x"18", x"18", x"18",
        x"00", x"00", x"00", x"00", x"38", x"44", x"44", x"44", x"38", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"78", x"44", x"44", x"44", x"78", x"40", x"40", x"00", x"00", x"08", x"10", x"20",
        x"00", x"00", x"00", x"00", x"3c", x"44", x"44", x"44", x"3c", x"04", x"04", x"00", x"20", x"20", x"10", x"08",
        x"00", x"00", x"00", x"00", x"58", x"64", x"40", x"40", x"40", x"00", x"00", x"00", x"00", x"08", x"04", x"02",
        x"00", x"00", x"00", x"00", x"3c", x"40", x"38", x"04", x"78", x"00", x"00", x"00", x"02", x"02", x"04", x"08",
        x"00", x"00", x"20", x"20", x"70", x"20", x"20", x"24", x"18", x"00", x"00", x"00", x"00", x"00", x"08", x"1C",
        x"00", x"00", x"00", x"00", x"44", x"44", x"44", x"4c", x"34", x"00", x"00", x"00", x"3E", x"1C", x"08", x"00",
        x"00", x"00", x"00", x"00", x"44", x"44", x"44", x"28", x"10", x"00", x"00", x"00", x"00", x"00", x"08", x"08",
        x"00", x"00", x"00", x"00", x"44", x"54", x"54", x"28", x"28", x"00", x"00", x"00", x"3E", x"08", x"08", x"00",
        x"00", x"00", x"00", x"00", x"44", x"28", x"10", x"28", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"00", x"00", x"44", x"44", x"44", x"3c", x"04", x"38", x"00", x"00", x"30", x"30", x"10", x"20",
        x"00", x"00", x"00", x"00", x"7c", x"08", x"10", x"20", x"7c", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"08", x"10", x"10", x"20", x"10", x"10", x"08", x"00", x"00", x"00", x"3E", x"00", x"00", x"00",
        x"00", x"00", x"10", x"10", x"10", x"00", x"10", x"10", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
        x"00", x"00", x"20", x"10", x"10", x"08", x"10", x"10", x"20", x"00", x"00", x"00", x"00", x"00", x"30", x"30",
        x"00", x"00", x"20", x"54", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"02", x"02", x"04",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"7c", x"00", x"00", x"00", x"08", x"10", x"20", x"20",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"24", x"24",
        x"00", x"00", x"00", x"08", x"00", x"08", x"08", x"08", x"08", x"08", x"00", x"00", x"24", x"24", x"24", x"18",
        x"00", x"00", x"00", x"00", x"08", x"1c", x"20", x"20", x"20", x"1c", x"08", x"00", x"00", x"08", x"18", x"08",
        x"00", x"00", x"00", x"0c", x"12", x"10", x"38", x"10", x"10", x"3e", x"00", x"00", x"08", x"08", x"08", x"1C",
        x"00", x"00", x"00", x"00", x"00", x"22", x"1c", x"14", x"1c", x"22", x"00", x"00", x"00", x"1C", x"22", x"02",
        x"00", x"00", x"00", x"22", x"14", x"08", x"3e", x"08", x"3e", x"08", x"00", x"00", x"1C", x"20", x"20", x"3E",
        x"00", x"00", x"00", x"08", x"08", x"08", x"00", x"08", x"08", x"08", x"00", x"00", x"00", x"1C", x"22", x"02",
        x"00", x"00", x"00", x"1c", x"20", x"1c", x"22", x"1c", x"02", x"1c", x"00", x"00", x"04", x"02", x"22", x"1C",
        x"14", x"14", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"14",
        x"00", x"00", x"3e", x"41", x"5d", x"51", x"51", x"5d", x"41", x"3e", x"00", x"00", x"3E", x"04", x"04", x"04",
        x"00", x"00", x"00", x"1c", x"02", x"1e", x"22", x"1e", x"00", x"00", x"00", x"00", x"00", x"3E", x"20", x"3C",
        x"00", x"00", x"00", x"00", x"0a", x"14", x"28", x"14", x"0a", x"00", x"00", x"00", x"02", x"02", x"22", x"1C",
        x"00", x"00", x"00", x"00", x"00", x"00", x"3e", x"02", x"02", x"00", x"00", x"00", x"00", x"1C", x"20", x"20",
        x"00", x"00", x"00", x"00", x"00", x"00", x"3e", x"00", x"00", x"00", x"00", x"00", x"3C", x"22", x"22", x"1C",
        x"00", x"00", x"3e", x"41", x"5d", x"55", x"59", x"55", x"41", x"3e", x"00", x"00", x"00", x"3E", x"02", x"04",
        x"00", x"00", x"00", x"7e", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"10", x"20", x"20",
        x"00", x"00", x"00", x"10", x"28", x"10", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"1C", x"22", x"22",
        x"00", x"00", x"08", x"08", x"3e", x"08", x"08", x"00", x"3e", x"00", x"00", x"00", x"1C", x"22", x"22", x"1C",
        x"00", x"00", x"00", x"18", x"04", x"08", x"10", x"1c", x"00", x"00", x"00", x"00", x"00", x"1C", x"22", x"22",
        x"00", x"00", x"00", x"18", x"04", x"18", x"04", x"18", x"00", x"00", x"00", x"00", x"1E", x"02", x"02", x"1C",
        x"04", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18",
        x"00", x"00", x"00", x"00", x"00", x"12", x"12", x"12", x"12", x"1c", x"10", x"20", x"00", x"18", x"18", x"00",
        x"00", x"00", x"00", x"1a", x"2a", x"2a", x"1a", x"0a", x"0a", x"0a", x"00", x"00", x"00", x"18", x"18", x"00",
        x"00", x"00", x"00", x"00", x"00", x"00", x"18", x"18", x"00", x"00", x"00", x"00", x"18", x"18", x"08", x"10",
        x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"18", x"00", x"04", x"08", x"10",
        x"00", x"00", x"00", x"08", x"18", x"08", x"08", x"1c", x"00", x"00", x"00", x"00", x"20", x"10", x"08", x"04",
        x"00", x"00", x"00", x"1c", x"22", x"22", x"22", x"1c", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"3E",
        x"00", x"00", x"00", x"00", x"28", x"14", x"0a", x"14", x"28", x"00", x"00", x"00", x"00", x"3E", x"00", x"00",
        x"00", x"00", x"00", x"20", x"20", x"20", x"22", x"06", x"0e", x"02", x"00", x"00", x"00", x"10", x"08", x"04",
        x"00", x"00", x"00", x"20", x"20", x"20", x"2e", x"02", x"04", x"0e", x"00", x"00", x"02", x"04", x"08", x"10",
        x"00", x"00", x"00", x"70", x"10", x"70", x"12", x"76", x"0e", x"02", x"00", x"00", x"00", x"18", x"24", x"04",
        x"00", x"00", x"00", x"08", x"00", x"08", x"08", x"10", x"12", x"0c", x"00", x"00", x"08", x"08", x"00", x"08"
    );

--attribute RAM_STYLE : string;
--attribute RAM_STYLE of RAM: signal is "BLOCK";

begin

    process (clka)
    begin
        if rising_edge(clka) then
            if (wea = '1') then
                RAM(conv_integer(addra(10 downto 0))) := dina;
            end if;
            douta <= RAM(conv_integer(addra(10 downto 0)));
        end if;
    end process;

    process (clkb)
    begin
        if rising_edge(clkb) then
            if (web = '1') then
                RAM(conv_integer(addrb(10 downto 0))) := dinb;
            end if;
            doutb <= RAM(conv_integer(addrb(10 downto 0)));
        end if;
    end process;

end BEHAVIORAL;

